module font_bitmap( input [3:0] x,
					input [3:0] y,
					input [3:0] digit,
					output pixel);
		
	wire[15:0] pattern;
	assign pixel = pattern[~x];
	
	assign pattern = 
		(digit == 4'd0) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000000000000
				:(y == 4'd2) ? 16'b0000111111100000
				:(y == 4'd3) ? 16'b0001110011110000
				:(y == 4'd4) ? 16'b0011100000111000
				:(y == 4'd5) ? 16'b0011000000011000
				:(y == 4'd6) ? 16'b0111000000011100
				:(y == 4'd7) ? 16'b0111000000011100
				:(y == 4'd8) ? 16'b0111000000111100
				:(y == 4'd9) ? 16'b0111000000111100
				:(y == 4'd10) ? 16'b0111100000111000
				:(y == 4'd11) ? 16'b0111111001111000
				:(y == 4'd12) ? 16'b0011111111111000
				:(y == 4'd13) ? 16'b0000111111110000
				:(y == 4'd14) ? 16'b0000001111000000
				: 16'b0000000000000000
				)
		:(digit == 4'd1) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0001000000000000
				:(y == 4'd2) ? 16'b0011111110000000
				:(y == 4'd3) ? 16'b0000000110000000
				:(y == 4'd4) ? 16'b0000000110000000
				:(y == 4'd5) ? 16'b0000000110000000
				:(y == 4'd6) ? 16'b0000000110000000
				:(y == 4'd7) ? 16'b0000000110000000
				:(y == 4'd8) ? 16'b0000001110000000
				:(y == 4'd9) ? 16'b0000001110000000
				:(y == 4'd10) ? 16'b0000001110000000
				:(y == 4'd11) ? 16'b0000001110000000
				:(y == 4'd12) ? 16'b0001111111111000
				:(y == 4'd13) ? 16'b0011111111111000
				:(y == 4'd14) ? 16'b0000000000000000
				:16'b0000000000000000
				)
		:(digit == 4'd2) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000000000000
				:(y == 4'd2) ? 16'b0000111111100000
				:(y == 4'd3) ? 16'b0001100000111000
				:(y == 4'd4) ? 16'b0011000000011000
				:(y == 4'd5) ? 16'b0011000000011000
				:(y == 4'd6) ? 16'b0000000000111000
				:(y == 4'd7) ? 16'b0000000001110000
				:(y == 4'd8) ? 16'b0000000111100000
				:(y == 4'd9) ? 16'b0000011100000000
				:(y == 4'd10) ? 16'b0001110000000000
				:(y == 4'd11) ? 16'b0011100000000000
				:(y == 4'd12) ? 16'b0011111111111000
				:(y == 4'd13) ? 16'b0011111111111000
				:(y == 4'd14) ? 16'b0000000000000000
				:16'b0000000000000000
				)
		:(digit == 4'd3) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000000000000
				:(y == 4'd2) ? 16'b0001111111111000
				:(y == 4'd3) ? 16'b0011111111110000
				:(y == 4'd4) ? 16'b0000000001100000
				:(y == 4'd5) ? 16'b0000000111000000
				:(y == 4'd6) ? 16'b0000001110000000
				:(y == 4'd7) ? 16'b0000011101110000
				:(y == 4'd8) ? 16'b0000010000011000
				:(y == 4'd9) ? 16'b0000000000011000
				:(y == 4'd10) ? 16'b0000000000011000
				:(y == 4'd11) ? 16'b0000000000111000
				:(y == 4'd12) ? 16'b0000000001110000
				:(y == 4'd13) ? 16'b0000000111100000
				:(y == 4'd14) ? 16'b0000111111000000
				: 16'b0001111100000000
				)
		:(digit == 4'd4) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000011000000
				:(y == 4'd2) ? 16'b0000000111000000
				:(y == 4'd3) ? 16'b0000000111000000
				:(y == 4'd4) ? 16'b0000001011000000
				:(y == 4'd5) ? 16'b0000011011000000
				:(y == 4'd6) ? 16'b0000110011000000
				:(y == 4'd7) ? 16'b0001110011000000
				:(y == 4'd8) ? 16'b0001100011000000
				:(y == 4'd9) ? 16'b0011111111100000
				:(y == 4'd10) ? 16'b0011111111111000
				:(y == 4'd11) ? 16'b0000000011100000
				:(y == 4'd12) ? 16'b0000000011000000
				:(y == 4'd13) ? 16'b0000000011000000
				:(y == 4'd14) ? 16'b0000000011000000
				: 16'b0000000000000000
				)
		:(digit == 4'd5) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0001111111111000
				:(y == 4'd2) ? 16'b0001111000000000
				:(y == 4'd3) ? 16'b0001100000000000
				:(y == 4'd4) ? 16'b0001100000000000
				:(y == 4'd5) ? 16'b0001111111100000
				:(y == 4'd6) ? 16'b0001111001110000
				:(y == 4'd7) ? 16'b0000000000011000
				:(y == 4'd8) ? 16'b0000000000011000
				:(y == 4'd9) ? 16'b0000000000011000
				:(y == 4'd10) ? 16'b0000000000110000
				:(y == 4'd11) ? 16'b0000000001100000
				:(y == 4'd12) ? 16'b0000001111000000
				:(y == 4'd13) ? 16'b0001111110000000
				:(y == 4'd14) ? 16'b0001110000000000
				: 16'b0000000000000000
				)
		:(digit == 4'd6) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000111110000
				:(y == 4'd2) ? 16'b0000011111110000
				:(y == 4'd3) ? 16'b0000111000000000
				:(y == 4'd4) ? 16'b0001110000000000
				:(y == 4'd5) ? 16'b0001100000000000
				:(y == 4'd6) ? 16'b0011001110000000
				:(y == 4'd7) ? 16'b0011111111100000
				:(y == 4'd8) ? 16'b0011100000110000
				:(y == 4'd9) ? 16'b0011000000010000
				:(y == 4'd10) ? 16'b0011000000011000
				:(y == 4'd11) ? 16'b0011000000011000
				:(y == 4'd12) ? 16'b0001110001110000
				:(y == 4'd13) ? 16'b0000111111100000
				:(y == 4'd14) ? 16'b0000000000000000
				: 16'b0000000000000000
				)
		:(digit == 4'd7) ? (
				(y == 4'd0) ? 16'b0011111111111000
				:(y == 4'd1) ? 16'b0011111111111000
				:(y == 4'd2) ? 16'b0011000000111000
				:(y == 4'd3) ? 16'b0010000001110000
				:(y == 4'd4) ? 16'b0000000001100000
				:(y == 4'd5) ? 16'b0000000011000000
				:(y == 4'd6) ? 16'b0000000011000000
				:(y == 4'd7) ? 16'b0000000110000000
				:(y == 4'd8) ? 16'b0000000110000000
				:(y == 4'd9) ? 16'b0000001110000000
				:(y == 4'd10) ? 16'b0000001110000000
				:(y == 4'd11) ? 16'b0000001110000000
				:(y == 4'd12) ? 16'b0000001100000000
				:(y == 4'd13) ? 16'b0000001100000000
				:(y == 4'd14) ? 16'b0000001100000000
				: 16'b0000000000000000
				)
		:(digit == 4'd8) ? (
				(y == 4'd0) ? 16'b0000001100000000
				:(y == 4'd1) ? 16'b0000111111100000
				:(y == 4'd2) ? 16'b0001110000110000
				:(y == 4'd3) ? 16'b0001100000011000
				:(y == 4'd4) ? 16'b0001100000011000
				:(y == 4'd5) ? 16'b0000110000110000
				:(y == 4'd6) ? 16'b0000111111110000
				:(y == 4'd7) ? 16'b0001111111110000
				:(y == 4'd8) ? 16'b0011100000011000
				:(y == 4'd9) ? 16'b0011000000001000
				:(y == 4'd10) ? 16'b0011000000001100
				:(y == 4'd11) ? 16'b0011000000011100
				:(y == 4'd12) ? 16'b0001110000111000
				:(y == 4'd13) ? 16'b0001111111110000
				:(y == 4'd14) ? 16'b0000001110000000
				: 16'b0000000000000000
				)
		:(digit == 4'd9) ? (
				(y == 4'd0) ? 16'b0000001110000000
				:(y == 4'd1) ? 16'b0000111111100000
				:(y == 4'd2) ? 16'b0001110011110000
				:(y == 4'd3) ? 16'b0011000000111000
				:(y == 4'd4) ? 16'b0011000000011000
				:(y == 4'd5) ? 16'b0011000000011000
				:(y == 4'd6) ? 16'b0011100000111000
				:(y == 4'd7) ? 16'b0001111111111000
				:(y == 4'd8) ? 16'b0000111111011000
				:(y == 4'd9) ? 16'b0000000000011000
				:(y == 4'd10) ? 16'b0000000000010000
				:(y == 4'd11) ? 16'b0000000000110000
				:(y == 4'd12) ? 16'b0000000011100000
				:(y == 4'd13) ? 16'b0001111111000000
				:(y == 4'd14) ? 16'b0001111000000000
				:16'b0000000000000000
				)
		:(digit == 4'd10) ? (
				(y == 4'd0) ?   16'b0000000000000000
				:(y == 4'd1) ?  16'b0000000000000000
				:(y == 4'd2) ?  16'b0000000000000000
				:(y == 4'd3) ?  16'b0000000000000000
				:(y == 4'd4) ?  16'b0000000100000000
				:(y == 4'd5) ?  16'b0000001110000000
				:(y == 4'd6) ?  16'b0000011011000000
				:(y == 4'd7) ?  16'b0000110001000000
				:(y == 4'd8) ?  16'b0000110001100000
				:(y == 4'd9) ?  16'b0000110001100000
				:(y == 4'd10) ? 16'b0000111111100000
				:(y == 4'd11) ? 16'b0001100001110000
				:(y == 4'd12) ? 16'b0111110000110000
				:(y == 4'd13) ? 16'b1111110011111110
				:(y == 4'd14) ? 16'b0000000000000000
				: 16'b0000000000000000
				)
		:(digit == 4'd11) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000000000000
				:(y == 4'd2) ? 16'b0111111111100000
				:(y == 4'd3) ? 16'b0111111111111000
				:(y == 4'd4) ? 16'b0000110000011000
				:(y == 4'd5) ? 16'b0000110000011000
				:(y == 4'd6) ? 16'b0000110000011000
				:(y == 4'd7) ? 16'b00001110111110000
				:(y == 4'd8) ? 16'b0000110000111000
				:(y == 4'd9) ? 16'b0000110000001100
				:(y == 4'd10) ? 16'b0000110000001100
				:(y == 4'd11) ? 16'b0000110000001100
				:(y == 4'd12) ? 16'b0000111111111000
				:(y == 4'd13) ? 16'b0111111111110000
				:(y == 4'd14) ? 16'b0000000000000000
				: 16'b0000000000000000
				)
		:(digit == 4'd12) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000000000000
				:(y == 4'd2) ? 16'b0000011111111000
				:(y == 4'd3) ? 16'b0000111001111000
				:(y == 4'd4) ? 16'b0001100000011000
				:(y == 4'd5) ? 16'b0011000000011000
				:(y == 4'd6) ? 16'b0011000000011000
				:(y == 4'd7) ? 16'b0011000000000000
				:(y == 4'd8) ? 16'b0011000000000000
				:(y == 4'd9) ? 16'b0011000000001000
				:(y == 4'd10) ? 16'b0001100000011000
				:(y == 4'd11) ? 16'b0001100000111000
				:(y == 4'd12) ? 16'b0000111111111000
				:(y == 4'd13) ? 16'b0000011111100000
				:(y == 4'd14) ? 16'b0000000000000000
				: 16'b0000000000000000
				)
		:(digit == 4'd13) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000000000000
				:(y == 4'd2) ? 16'b0111111111100000
				:(y == 4'd3) ? 16'b0000111000110000
				:(y == 4'd4) ? 16'b0000110000011000
				:(y == 4'd5) ? 16'b0000110000001100
				:(y == 4'd6) ? 16'b0000110000000110
				:(y == 4'd7) ? 16'b0000110000000110
				:(y == 4'd8) ? 16'b0000110000000110
				:(y == 4'd9) ? 16'b0000110000000110
				:(y == 4'd10) ? 16'b0000110000001100
				:(y == 4'd11) ? 16'b0000110000001100
				:(y == 4'd12) ? 16'b0000110000111000
				:(y == 4'd13) ? 16'b0111111111100000
				:(y == 4'd14) ? 16'b0010000000000000
				: 16'b0000000000000000
				)
		:(digit == 4'd14) ? (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000000000000
				:(y == 4'd2) ? 16'b0111111111111000
				:(y == 4'd3) ? 16'b0000110000001100
				:(y == 4'd4) ? 16'b0000110000000100
				:(y == 4'd5) ? 16'b0000110001100100
				:(y == 4'd6) ? 16'b0000110011100000
				:(y == 4'd7) ? 16'b0000111111100000
				:(y == 4'd8) ? 16'b0000110001100000
				:(y == 4'd9) ? 16'b0000110001000100
				:(y == 4'd10) ? 16'b0000110000000110
				:(y == 4'd11) ? 16'b0000110000001100
				:(y == 4'd12) ? 16'b0011111111111100
				:(y == 4'd13) ? 16'b0111111111111100
				:(y == 4'd14) ? 16'b0000000000000000
				: 16'b0000000000000000
				)
		: (
				(y == 4'd0) ? 16'b0000000000000000
				:(y == 4'd1) ? 16'b0000000000000000
				:(y == 4'd2) ? 16'b0011111111110000
				:(y == 4'd3) ? 16'b0111111111111100
				:(y == 4'd4) ? 16'b0000110000001110
				:(y == 4'd5) ? 16'b0000110000000100
				:(y == 4'd6) ? 16'b0000110001000000
				:(y == 4'd7) ? 16'b0000111111000000
				:(y == 4'd8) ? 16'b0000111100000000
				:(y == 4'd9) ? 16'b0000110000000000
				:(y == 4'd10) ? 16'b0000110000000000
				:(y == 4'd11) ? 16'b0000110000000000
				:(y == 4'd12) ? 16'b0000110000000000
				:(y == 4'd13) ? 16'b0011111111000000
				:(y == 4'd14) ? 16'b0010000000000000
				: 16'b0000000000000000
				);
endmodule