module myrom(input clk, input[4:0] addr, output reg [439:0] data);
always @(posedge clk) 
case (addr)
	5'd0 : data <= 440'h 45F7612A1CEC52E70385A02EF721FCFAA3DC18B1EFF7E89BF76786329C4813DFA3276C941F3680745FAAB1F6F4414F427E1D6FD7EF98F8;
	5'd1 : data <= 440'h 13F9A11ABADBD605D355E8CDC8D93D4A88B3E558EF7612F6694CE752B67A4ED025BB38965D2AA9AEB5E299DB3872F8E55D1D766473B336;
	5'd2 : data <= 440'h A6EEDE6FB39CD2988855324137380692AB48F9EF732F5C3FA212B90528B0CB1F40EA63B3FB206B828019B0684C791102523A63F1369E52;
	5'd3 : data <= 440'h 9896C52DD1FE93304F41BAE8245D5D283E49377820195C8E67781B68F3E9433B9C344AB890F8D2C17BA35D2742074D1330B02FECC3AB96;
	5'd4 : data <= 440'h A5505C3AE01A164FC35D905429B427E646421B28E9E0E2ACA462573821E16064E642FFB3198E168D6755C536746FFE31F3676489DC4F7C;
	5'd5 : data <= 440'h 2DBB48CC248E266AB90E83F490C043F29A331B76F8ECE93E7E313EC7F870D460EDA886D9ECC196EA3765FBC2CD6A4339650340C79E0B8F;
	5'd6 : data <= 440'h 29B6C18975D92E49E90FF9E211002870D2C92C87003FCFF55CCBA1D5E7C5FCE4D0FE89160EFF8EDEFD6A854AB42E6F5870A94BAD96EE16;
	5'd7 : data <= 440'h 58220D18D3AB86398316E646E7E05723DB3FE533FF94C12502B145C9D47124BC9CB12576FB84745AA1927848770571CCE1039C0C94579C;
	5'd8 : data <= 440'h 5BCFE0779BD58963DA4D56E4C84527FC1C72A98F7733050AE2A4BD80CAF5422EE3E4517542397DCE764595B17FF677EA08C6DA0993C865;
	5'd9 : data <= 440'h 310C5BAB3CC04B1DF9BEFF6D2F9C0D092C59D2F895F783FAB56A353366FEECD4627B212C241D53DB49A5D380DF8CEB8E70AB1FECEFFC95;
	5'd10 : data <= 440'h 1502A9DCD6E64FC5FD5420F2BADA828532A453289BD47B363738F8662D2C6EED07CB8B892FCE0F4832D99AAA20B2B82FD1E1355E442CBA;
	5'd11 : data <= 440'h 4162A7A77D6957FA7BB3345BF595EB8A8FC7C1F2A46626CF17C40BC6888C4C8234A03BBF0B5AACA2BD81E430F65FB4FACEAF8D2542F07D;
	5'd12 : data <= 440'h 8432ECC0D215B5BD1B7B2533E19A99A8B404DA6FEABE3A3B4A5426376B55BAC3744A6B50E5C68238E582BBC62199ACC30A932B7EB65BAA;
	5'd13 : data <= 440'h 7A0FC160C9DA40940C964642A9EC0B9BC2929F2A2A38C9D003AE5B45D32BFC4C154893705BEAD78E54059A17CB4FAFF9A9F0C04F81E0A2;
	5'd14 : data <= 440'h 58CC28DD5DB9408728BF4BC92CC4D50B638D8454A6854741126C4A01B3023D7D7330CB3E4E5DDC66168CEACF59BA6D2DAC1861723F5C7D;
	5'd15 : data <= 440'h 390EE7B13A7C99B739227452AA30B9864B7A4C83290855C8FFC55BC3C0BCA532B832881E4B945728D1244303D272BF7E7B0E1EEF140475;
	5'd16 : data <= 440'h 53C78DED178A72C15BBF3451248922DD36A9965916287D08D8E2ECE048980AAE3175E0073E9B6E7E615302B6FDE42FF660BF14890380A6;
	5'd17 : data <= 440'h 8D9359D087CA6E6B870B97C5E1C97363204E5335E697F7398A9ECEB219EDCDB25D46600666C6DE66C5E9298C6C44EAF02BD18A15AFAF25;
	5'd18 : data <= 440'h 8E6E244EA54621021773C8BCBEC24198B0C3207D3458A2E1539A16F03F26CAA2196AE32D294CE78BF3657C141A42CBC5C4DE8086F8F80F;
	5'd19 : data <= 440'h 1460922C2AC80434C9828D117D69D1899B8E544F05C6DE4756B8B09280B3D49580BAE10A4972770C9D5C650A82C33F0C89C80E8A5D4360;
	5'd20 : data <= 440'h 3A9FD5EAAC281AE234ACC416E55C4EC7172C76B92D315D164F26C0488E44824FC16504AB169F3821A8A437B98EDB8FFE4A73E3FD75BEDD;
	5'd21 : data <= 440'h 96B6FA91EFAB3A16277426F6620800094AE3410622CD598ED3E74AB9B6FE34B50EEC605FB384D9E0AF1C719A45FC7566E29FC0D5AE37AE;
	5'd22 : data <= 440'h 3B6EF3202C602060BD7ABADDDCD4061CE46D6DF12EC86F376377B518EE20863C8D101452AE09C77B63DA12C25EA761EBE3A678D88387D1;
	5'd23 : data <= 440'h 9022F0D689BDA25E1D6C884EB1A93273F5EC1A26FCC9D7DF3C448F45F8E510DFF1060A570B2F4EB79D068B501FE09E0406557E8BE04355;
	5'd24 : data <= 440'h 812D5307CC9301CC207CE0E01C64C84A14EBEF82079FF92946188EB15B73E0B1186961592AF6D1B81C881EE1942BAA03AE811AF8EBAD5D;
	5'd25 : data <= 440'h 9A77C9F992FE656809ADC7FD8C752B0B83BE497F42B1776C84ACD0E5E0E43C9E2E875A62A74A251BA58C4C60540311A59113E00262EF24;
	5'd26 : data <= 440'h 952ADB04CD26E59C71EEF394E2055BB500D476FAB7A907CB7D58884AC04CB36E41FDF4BDF944A3450E60B308E198AF763B76DBB7DF6309;
	5'd27 : data <= 440'h B63BF394566ED3E5A44DD20DC884AE694E55595D939AA4522BF69970793A7E877F1D2CDCED81C624441816FFB7B7F9C5855901BA901EF;
	5'd28 : data <= 440'h 2B12A18F32819A5CBE8C87A061D0A71054A857FB1034B61DA0412B95C1487DD0CBF3BC93F1CFA3D70F18500EAE0BBD684CEA9D621429B6;
	5'd29 : data <= 440'h 7A40B4F057560B111B67A4BBB2D66B69D7EB5C50BC8C63238B615EB158867EE9C1307B463D91AE745B0A5BAEACD006F24DC9BABB74D92B;
	5'd30 : data <= 440'h 898C6989448FAFA73C2E30509191817EAE0633B99B178EC507DFCE60B45177CC7F574483FA2B4F60ECA6F34B5B9331370ABE66ECE0DFF8;
	5'd31 : data <= 440'h C9467949D89A9FA9CD6D5166D9051B36BD6547B986B04B55ADBD04A478C54E31FF41AC2005ABD3AAD03C8CB2109CC05981D227D013FEE;
endcase
endmodule

module Randomwalk_ROM(input clk, input[7:0] addr, output reg [109:0] data);
always @(posedge clk)
	case (addr)
		8'd0	: data	<= 110'h11174AE60A7E8B7C46574CE4FDFF;
		8'd1	: data	<= 110'h0;
		8'd2	: data	<= 110'hC72AD1A1D30AF27B057AB643BBC;
		8'd3	: data	<= 110'h7B1992EABF13F43CEC85203222D;
		8'd4	: data	<= 110'h2;
		8'd5	: data	<= 110'h0;
		8'd6	: data	<= 110'h12782F269E06F34D7BB4F4E5645B;
		8'd7	: data	<= 110'h1EBFC2FC5154F1EF61A488B44DF3;
		8'd8	: data	<= 110'h4;
		8'd9	: data	<= 110'h0;
		8'd10	: data	<= 110'hA9C209480C1E1808D6E80F6E143;
		8'd11	: data	<= 110'h1A98F92699F796384B7EAB43242;
		8'd12	: data	<= 110'h8;
		8'd13	: data	<= 110'h0;
		8'd14	: data	<= 110'h68C48C85B8E02D3F781B67554D2;
		8'd15	: data	<= 110'hB4708162617FA04349DBB47D89E;
		8'd16	: data	<= 110'h10;
		8'd17	: data	<= 110'h0;
		8'd18	: data	<= 110'h23A850E12934537B74AC50CFF407;
		8'd19	: data	<= 110'h8B427B17A481C1270550E2C9795;
		8'd20	: data	<= 110'h20;
		8'd21	: data	<= 110'h0;
		8'd22	: data	<= 110'h2BA31DEEBA75F0AA2E193A5B4A4F;
		8'd23	: data	<= 110'h12879B85F258ED2274ED70A9F172;
		8'd24	: data	<= 110'h40;
		8'd25	: data	<= 110'h0;
		8'd26	: data	<= 110'h253EE2BC8E247CF8E9B762E7D2B4;
		8'd27	: data	<= 110'h2D9DC156B7A376EB6DF35590628;
		8'd28	: data	<= 110'h80;
		8'd29	: data	<= 110'h0;
		8'd30	: data	<= 110'h1E69227CBE1F7616DDE2A33ADD83;
		8'd31	: data	<= 110'h26C828150B1D30F0D7B0F5C70A46;
		8'd32	: data	<= 110'h100;
		8'd33	: data	<= 110'h0;
		8'd34	: data	<= 110'h14C29315BDECDF18DC31D0F5E407;
		8'd35	: data	<= 110'h1A466B668B1ED335EE1CABA73BA8;
		8'd36	: data	<= 110'h200;
		8'd37	: data	<= 110'h0;
		8'd38	: data	<= 110'h271230736F199B011A413C156CF1;
		8'd39	: data	<= 110'h2365F19901AAF99595632F6EDD72;
		8'd40	: data	<= 110'h400;
		8'd41	: data	<= 110'h0;
		8'd42	: data	<= 110'h7D62EEE76DE1D904E7723AB74C3;
		8'd43	: data	<= 110'hA67452070B9122F4AB3387AB51B;
		8'd44	: data	<= 110'h800;
		8'd45	: data	<= 110'h0;
		8'd46	: data	<= 110'h94C0A3FEDDB5A67589C168EFB18;
		8'd47	: data	<= 110'h117D9822ED6D0EC1D6CC32A12F1F;
		8'd48	: data	<= 110'h1000;
		8'd49	: data	<= 110'h0;
		8'd50	: data	<= 110'h15546F88615CA582BFFDE4E7BDB;
		8'd51	: data	<= 110'hBC6B6703075890A4A7AB32404FC;
		8'd52	: data	<= 110'h2000;
		8'd53	: data	<= 110'h0;
		8'd54	: data	<= 110'h56FC974556EDE3A32BEA9D7A1A8;
		8'd55	: data	<= 110'h47B8F2B5E717894644BAFB9653C;
		8'd56	: data	<= 110'h4000;
		8'd57	: data	<= 110'h0;
		8'd58	: data	<= 110'h10C3A9D7DABDD18D28ADC6FB94E3;
		8'd59	: data	<= 110'hE4772AB18C0F1EB697BE9693740;
		8'd60	: data	<= 110'h8000;
		8'd61	: data	<= 110'h0;
		8'd62	: data	<= 110'hDAA83A0032095CB94E36F89D3B8;
		8'd63	: data	<= 110'hD80BBEF77CE7C5068425DF1E5DE;
		8'd64	: data	<= 110'h10000;
		8'd65	: data	<= 110'h0;
		8'd66	: data	<= 110'h244F12D3F1BFE534A9BB5BE9B823;
		8'd67	: data	<= 110'h2B3691F6B73E90C84ECC1A14FF1E;
		8'd68	: data	<= 110'h20000;
		8'd69	: data	<= 110'h0;
		8'd70	: data	<= 110'h24C54FC5E8569AE8EFD8F2EAC4D9;
		8'd71	: data	<= 110'h2037CB37D60C96543B7D3C9C7CCB;
		8'd72	: data	<= 110'h40000;
		8'd73	: data	<= 110'h0;
		8'd74	: data	<= 110'h1CBAF3CE0FD34583F329401F0C5;
		8'd75	: data	<= 110'h2645B1D2DD72547B11A30CE8B3FD;
		8'd76	: data	<= 110'h80000;
		8'd77	: data	<= 110'h0;
		8'd78	: data	<= 110'h3C76BB97F733B825AF36B1DB980;
		8'd79	: data	<= 110'h1CE7F1D1FA8F79AB74B7EFCBEAE3;
		8'd80	: data	<= 110'h100000;
		8'd81	: data	<= 110'h0;
		8'd82	: data	<= 110'h77FF7CFB5EE44C62072CFD09A21;
		8'd83	: data	<= 110'h20AF72D276437457EEAB3FAC8C3B;
		8'd84	: data	<= 110'h200000;
		8'd85	: data	<= 110'h0;
		8'd86	: data	<= 110'h73DA67110FEE3BE369565B718A2;
		8'd87	: data	<= 110'h94DAC4C858CE1D1676C9CFAF526;
		8'd88	: data	<= 110'h400000;
		8'd89	: data	<= 110'h0;
		8'd90	: data	<= 110'h17F84CE7E8B3882A89823DD40540;
		8'd91	: data	<= 110'h26ABAF7BCB98391B4C52E2139BA4;
		8'd92	: data	<= 110'h800000;
		8'd93	: data	<= 110'h0;
		8'd94	: data	<= 110'h25871DB9C2D7427EA6E84655A50F;
		8'd95	: data	<= 110'h288432D0DFF687FC2EB1A7B828B4;
		8'd96	: data	<= 110'h1000000;
		8'd97	: data	<= 110'h0;
		8'd98	: data	<= 110'h6CE7AF6674207ACD7BC21472BA7;
		8'd99	: data	<= 110'h15DCA7BA7937863AB3692545F6B8;
		8'd100	: data	<= 110'h2000000;
		8'd101	: data	<= 110'h0;
		8'd102	: data	<= 110'h511E6477C078315A6E0A5AC9233;
		8'd103	: data	<= 110'h20475274362CF41C9D4593B3AD40;
		8'd104	: data	<= 110'h4000000;
		8'd105	: data	<= 110'h0;
		8'd106	: data	<= 110'h719F7A8B5272B6495DDD6DBEE67;
		8'd107	: data	<= 110'h1F21BF0F8A0D5C66156BEEBAD344;
		8'd108	: data	<= 110'h8000000;
		8'd109	: data	<= 110'h0;
		8'd110	: data	<= 110'h171167D11502BC0034DDF16842A9;
		8'd111	: data	<= 110'h1F77A746567352996F6E0D150D01;
		8'd112	: data	<= 110'h10000000;
		8'd113	: data	<= 110'h0;
		8'd114	: data	<= 110'hBF96DA58A42BC03E8250A0B78F0;
		8'd115	: data	<= 110'h152038C4F62D7DD5E5707C0104CE;
		8'd116	: data	<= 110'h20000000;
		8'd117	: data	<= 110'h0;
		8'd118	: data	<= 110'h1BE903BEBD4FA1B629CBB6AB7C09;
		8'd119	: data	<= 110'hCC95694AA7F961F71B726F7A64;
		8'd120	: data	<= 110'h40000000;
		8'd121	: data	<= 110'h0;
		8'd122	: data	<= 110'h1623EA7EEE32BE90B37DD8D999D6;
		8'd123	: data	<= 110'hF46C132DA13D750BCC89DE1B5AD;
		8'd124	: data	<= 110'h80000000;
		8'd125	: data	<= 110'h0;
		8'd126	: data	<= 110'h26E28AFF1949A35B71DD3FFA6E38;
		8'd127	: data	<= 110'hCE0AB7C12530DB75008ECCE4D15;
		8'd128	: data	<= 110'h117DD84A873B14B9C0E1680BBDC8;
		8'd129	: data	<= 110'h1FCFAA3DC18B1EFF7E89BF767863;
		8'd130	: data	<= 110'hA71204F7E8C9DB2507CDA01D17E;
		8'd131	: data	<= 110'h2AB1F6F4414F427E1D6FD7EF98F8;
		8'd132	: data	<= 110'h4FE6846AEB6F58174D57A337236;
		8'd133	: data	<= 110'h13D4A88B3E558EF7612F6694CE75;
		8'd134	: data	<= 110'hAD9E93B4096ECE25974AAA6BAD7;
		8'd135	: data	<= 110'h2299DB3872F8E55D1D766473B336;
		8'd136	: data	<= 110'h29BBB79BECE734A622154C904DCE;
		8'd137	: data	<= 110'h692AB48F9EF732F5C3FA212B90;
		8'd138	: data	<= 110'h14A2C32C7D03A98ECFEC81AE0A00;
		8'd139	: data	<= 110'h19B0684C791102523A63F1369E52;
		8'd140	: data	<= 110'h2625B14B747FA4CC13D06EBA0917;
		8'd141	: data	<= 110'h15D283E49377820195C8E67781B6;
		8'd142	: data	<= 110'h23CFA50CEE70D12AE243E34B05EE;
		8'd143	: data	<= 110'h235D2742074D1330B02FECC3AB96;
		8'd144	: data	<= 110'h2954170EB8068593F0D764150A6D;
		8'd145	: data	<= 110'h27E646421B28E9E0E2ACA462573;
		8'd146	: data	<= 110'h2087858193990BFECC66385A359D;
		8'd147	: data	<= 110'h15C536746FFE31F3676489DC4F7C;
		8'd148	: data	<= 110'hB6ED2330923899AAE43A0FD2430;
		8'd149	: data	<= 110'h43F29A331B76F8ECE93E7E313EC;
		8'd150	: data	<= 110'h1FE1C35183B6A21B67B3065BA8DD;
		8'd151	: data	<= 110'h25FBC2CD6A4339650340C79E0B8F;
		8'd152	: data	<= 110'hA6DB0625D764B927A43FE788440;
		8'd153	: data	<= 110'h2870D2C92C87003FCFF55CCBA1D;
		8'd154	: data	<= 110'h179F17F39343FA24583BFE3B7BF5;
		8'd155	: data	<= 110'h2A854AB42E6F5870A94BAD96EE16;
		8'd156	: data	<= 110'h1608834634EAE18E60C5B991B9F8;
		8'd157	: data	<= 110'h5723DB3FE533FF94C12502B145C;
		8'd158	: data	<= 110'h2751C492F272C495DBEE11D16A86;
		8'd159	: data	<= 110'h127848770571CCE1039C0C94579C;
		8'd160	: data	<= 110'h16F3F81DE6F56258F69355B93211;
		8'd161	: data	<= 110'h127FC1C72A98F7733050AE2A4BD8;
		8'd162	: data	<= 110'h32BD508BB8F9145D508E5F739D9;
		8'd163	: data	<= 110'h595B17FF677EA08C6DA0993C865;
		8'd164	: data	<= 110'hC4316EACF3012C77E6FBFDB4BE7;
		8'd165	: data	<= 110'hD092C59D2F895F783FAB56A353;
		8'd166	: data	<= 110'hD9BFBB35189EC84B090754F6D26;
		8'd167	: data	<= 110'h25D380DF8CEB8E70AB1FECEFFC95;
		8'd168	: data	<= 110'h540AA7735B993F17F55083CAEB6;
		8'd169	: data	<= 110'h2828532A453289BD47B363738F86;
		8'd170	: data	<= 110'h18B4B1BBB41F2E2E24BF383D20CB;
		8'd171	: data	<= 110'h199AAA20B2B82FD1E1355E442CBA;
		8'd172	: data	<= 110'h1058A9E9DF5A55FE9EECCD16FD65;
		8'd173	: data	<= 110'h1EB8A8FC7C1F2A46626CF17C40BC;
		8'd174	: data	<= 110'h1A22313208D280EEFC2D6AB28AF6;
		8'd175	: data	<= 110'h1E430F65FB4FACEAF8D2542F07D;
		8'd176	: data	<= 110'h210CBB3034856D6F46DEC94CF866;
		8'd177	: data	<= 110'h299A8B404DA6FEABE3A3B4A54263;
		8'd178	: data	<= 110'h1DAD56EB0DD129AD43971A08E396;
		8'd179	: data	<= 110'h2BBC62199ACC30A932B7EB65BAA;
		8'd180	: data	<= 110'h1E83F0583276902503259190AA7B;
		8'd181	: data	<= 110'hB9BC2929F2A2A38C9D003AE5B4;
		8'd182	: data	<= 110'h174CAFF13055224DC16FAB5E3950;
		8'd183	: data	<= 110'h59A17CB4FAFF9A9F0C04F81E0A2;
		8'd184	: data	<= 110'h16330A37576E5021CA2FD2F24B31;
		8'd185	: data	<= 110'hD50B638D8454A6854741126C4A0;
		8'd186	: data	<= 110'h6CC08F5F5CCC32CF9397771985A;
		8'd187	: data	<= 110'hCEACF59BA6D2DAC1861723F5C7D;
		8'd188	: data	<= 110'hE43B9EC4E9F266DCE489D14AA8C;
		8'd189	: data	<= 110'hB9864B7A4C83290855C8FFC55BC;
		8'd190	: data	<= 110'hF02F294CAE0CA20792E515CA344;
		8'd191	: data	<= 110'h244303D272BF7E7B0E1EEF140475;
		8'd192	: data	<= 110'h14F1E37B45E29CB056EFCD144922;
		8'd193	: data	<= 110'h122DD36A9965916287D08D8E2ECE;
		8'd194	: data	<= 110'h122602AB8C5D7801CFA6DB9F985;
		8'd195	: data	<= 110'h1302B6FDE42FF660BF14890380A6;
		8'd196	: data	<= 110'h2364D67421F29B9AE1C2E5F17872;
		8'd197	: data	<= 110'h17363204E5335E697F7398A9ECEB;
		8'd198	: data	<= 110'h867B736C9751980199B1B799B17;
		8'd199	: data	<= 110'h29298C6C44EAF02BD18A15AFAF25;
		8'd200	: data	<= 110'h239B8913A951884085DCF22F2FB0;
		8'd201	: data	<= 110'h24198B0C3207D3458A2E1539A16F;
		8'd202	: data	<= 110'hFC9B2A8865AB8CB4A5339E2FCD;
		8'd203	: data	<= 110'h257C141A42CBC5C4DE8086F8F80F;
		8'd204	: data	<= 110'h518248B0AB2010D3260A3445F5A;
		8'd205	: data	<= 110'h1D1899B8E544F05C6DE4756B8B09;
		8'd206	: data	<= 110'hA02CF525602EB842925C9DC3275;
		8'd207	: data	<= 110'h1C650A82C33F0C89C80E8A5D4360;
		8'd208	: data	<= 110'hEA7F57AAB0A06B88D2B3105B957;
		8'd209	: data	<= 110'h4EC7172C76B92D315D164F26C04;
		8'd210	: data	<= 110'h223912093F059412AC5A7CE086A2;
		8'd211	: data	<= 110'h2437B98EDB8FFE4A73E3FD75BEDD;
		8'd212	: data	<= 110'h25ADBEA47BEACE8589DD09BD9882;
		8'd213	: data	<= 110'h94AE3410622CD598ED3E74AB;
		8'd214	: data	<= 110'h26DBF8D2D43BB1817ECE136782BC;
		8'd215	: data	<= 110'h1C719A45FC7566E29FC0D5AE37AE;
		8'd216	: data	<= 110'hEDBBCC80B1808182F5EAEB77735;
		8'd217	: data	<= 110'h61CE46D6DF12EC86F376377B51;
		8'd218	: data	<= 110'h23B88218F23440514AB8271DED8F;
		8'd219	: data	<= 110'h1A12C25EA761EBE3A678D88387D1;
		8'd220	: data	<= 110'h2408BC35A26F6897875B2213AC6A;
		8'd221	: data	<= 110'h13273F5EC1A26FCC9D7DF3C448F4;
		8'd222	: data	<= 110'h17E394437FC418295C2CBD3ADE74;
		8'd223	: data	<= 110'h68B501FE09E0406557E8BE04355;
		8'd224	: data	<= 110'h204B54C1F324C073081F38380719;
		8'd225	: data	<= 110'hC84A14EBEF82079FF92946188EB;
		8'd226	: data	<= 110'h56DCF82C461A58564ABDB46E072;
		8'd227	: data	<= 110'h81EE1942BAA03AE811AF8EBAD5D;
		8'd228	: data	<= 110'h269DF27E64BF995A026B71FF631D;
		8'd229	: data	<= 110'h12B0B83BE497F42B1776C84ACD0E;
		8'd230	: data	<= 110'h178390F278BA1D698A9D28946E96;
		8'd231	: data	<= 110'hC4C60540311A59113E00262EF24;
		8'd232	: data	<= 110'h254AB6C13349B9671C7BBCE53881;
		8'd233	: data	<= 110'h15BB500D476FAB7A907CB7D58884;
		8'd234	: data	<= 110'h2B0132CDB907F7D2F7E5128D1439;
		8'd235	: data	<= 110'h20B308E198AF763B76DBB7DF6309;
		8'd236	: data	<= 110'h2D8EFCE5159BB4F969137483722;
		8'd237	: data	<= 110'h4AE694E55595D939AA4522BF699;
		8'd238	: data	<= 110'h1C1E4E9FA1DFC74B373B60718911;
		8'd239	: data	<= 110'h1816FFB7B7F9C5855901BA901EF;
		8'd240	: data	<= 110'hAC4A863CCA066972FA321E81874;
		8'd241	: data	<= 110'hA71054A857FB1034B61DA0412B9;
		8'd242	: data	<= 110'h170521F7432FCEF24FC73E8F5C3C;
		8'd243	: data	<= 110'h18500EAE0BBD684CEA9D621429B6;
		8'd244	: data	<= 110'h1E902D3C15D582C446D9E92EECB5;
		8'd245	: data	<= 110'h26B69D7EB5C50BC8C63238B615EB;
		8'd246	: data	<= 110'h56219FBA704C1ED18F646B9D16C;
		8'd247	: data	<= 110'hA5BAEACD006F24DC9BABB74D92B;
		8'd248	: data	<= 110'h22631A625123EBE9CF0B8C142464;
		8'd249	: data	<= 110'h1817EAE0633B99B178EC507DFCE6;
		8'd250	: data	<= 110'h2D145DF31FD5D120FE8AD3D83B2;
		8'd251	: data	<= 110'h26F34B5B9331370ABE66ECE0DFF8;
		8'd252	: data	<= 110'h32519E527626A7EA735B5459B64;
		8'd253	: data	<= 110'h51B36BD6547B986B04B55ADBD04;
		8'd254	: data	<= 110'h291E31538C7FD06B08016AF4EAB4;
		8'd255	: data	<= 110'h3C8CB2109CC05981D227D013FEE;
	endcase
endmodule

